
module PiSimulator_VGA (
   
)
